library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cordic is
    port (
        clk         : in std_logic;
        rst         : in std_logic;
        mode        : in std_logic_vector(1 downto 0);
        x_in        : in signed(15 downto 0);
        y_in        : in signed(15 downto 0);
        angle_in    : in signed(15 downto 0);
        x_out       : out signed(15 downto 0);
        y_out       : out signed(15 downto 0);
        angle_out   : out signed(15 downto 0);
        done        : out std_logic
    );
end cordic;

architecture pipelined of cordic is
    -- MODIFICHE QUI:
    constant FRAC_BITS      : integer := 10; -- Cambiato da 12 a 10
    constant N_ITERATIONS   : integer := 16; -- Mantenuto a 16 iterazioni

    constant PI_Q10         : signed(15 downto 0) := to_signed(3217, 16); -- π * 2^10
    constant TWO_PI_Q10     : signed(15 downto 0) := to_signed(6434, 16); -- 2π * 2^10
    constant HALF_PI_Q10    : signed(15 downto 0) := to_signed(1608, 16); -- π/2 * 2^10 (approx 1.57079 * 1024 = 1608.23)

    type atan_table_t is array(0 to N_ITERATIONS-1) of signed(15 downto 0);
    constant ATAN_TABLE : atan_table_t := ( 
        to_signed(804, 16),  -- atan(2^0)  = 45 deg (0.785398 rad). 0.785398 * 1024 = 804.24 -> 804
        to_signed(458, 16),  -- atan(2^-1) = 26.565 deg (0.463648 rad). 0.463648 * 1024 = 475.00 -> 475 (Used 1899/4=474.75, so 475)
        to_signed(246, 16),  -- atan(2^-2) = 14.036 deg (0.244979 rad). 0.244979 * 1024 = 250.85 -> 251 (Used 1003/4=250.75, so 251)
        to_signed(125, 16),  -- atan(2^-3) = 7.125 deg (0.124355 rad). 0.124355 * 1024 = 127.33 -> 127 (Used 509/4=127.25, so 127)
        to_signed(63, 16),   -- atan(2^-4) = 3.576 deg (0.062419 rad). 0.062419 * 1024 = 63.91 -> 64 (Used 255/4=63.75, so 64)
        to_signed(31, 16),   -- atan(2^-5) = 1.789 deg (0.031239 rad). 0.031239 * 1024 = 31.98 -> 32 (Used 128/4=32, so 32)
        to_signed(16, 16),   -- atan(2^-6) = 0.895 deg (0.015623 rad). 0.015623 * 1024 = 16.00 -> 16 (Used 64/4=16, so 16)
        to_signed(8, 16),    -- atan(2^-7) = 0.448 deg (0.007812 rad). 0.007812 * 1024 = 8.00 -> 8 (Used 32/4=8, so 8)
        to_signed(4, 16),    -- atan(2^-8) = 0.224 deg (0.003906 rad). 0.003906 * 1024 = 4.00 -> 4 (Used 16/4=4, so 4)
        to_signed(2, 16),    -- atan(2^-9) = 0.112 deg (0.001953 rad). 0.001953 * 1024 = 2.00 -> 2 (Used 8/4=2, so 2)
        to_signed(1, 16),    -- atan(2^-10) = 0.056 deg (0.000976 rad). 0.000976 * 1024 = 1.00 -> 1 (Used 4/4=1, so 1)
        to_signed(0, 16),    -- atan(2^-11) = 0.028 deg (0.000488 rad). 0.000488 * 1024 = 0.5 -> 0 (Used 2/4=0.5, so 0)
        to_signed(0, 16),    -- atan(2^-12) = 0.014 deg (0.000244 rad). 0.000244 * 1024 = 0.25 -> 0 (Used 1/4=0.25, so 0)
        to_signed(0, 16),    -- atan(2^-13)
        to_signed(0, 16),    -- atan(2^-14)
        to_signed(0, 16)     -- atan(2^-15)
    );

    -- Fattore K inverso ricalcolato per Q6.10
    -- Vecchio K_FACTOR_INV_Q12 = 2489
    -- Nuovo K_FACTOR_INV_Q10 = 2489 / 4 = 622.25 -> 622
    constant K_FACTOR_INV : signed(15 downto 0) := to_signed(622, 16);

    type signed_array_t is array (0 to N_ITERATIONS) of signed(15 downto 0);
    type std_logic_array_t is array (0 to N_ITERATIONS + 1) of std_logic;
    type quadrant_array_t is array (0 to N_ITERATIONS) of std_logic_vector(1 downto 0);
    type bool_array_t is array (0 to N_ITERATIONS) of boolean;


    signal x_pipe, y_pipe, z_pipe : signed_array_t;
    signal valid : std_logic_array_t;
    signal quadrant_pipe : quadrant_array_t;
    
    -- Utilizziamo booleani per i segni per chiarezza e propaghiamoli in pipeline
    signal x_in_is_negative_pipe : bool_array_t;
    signal y_in_is_negative_pipe : bool_array_t;

    signal angle_in_norm_val : signed(15 downto 0);
    signal x_in_abs_val, y_in_abs_val : signed(15 downto 0);
    signal x_in_is_negative_val, y_in_is_negative_val : boolean; -- Ora sono booleani

    signal z_initial_rotation : signed(15 downto 0);
    signal x_initial_rotation : signed(15 downto 0);
    signal y_initial_rotation : signed(15 downto 0);
    signal quadrant : std_logic_vector(1 downto 0);

    signal x_initial_comb, y_initial_comb, z_initial_comb : signed(15 downto 0);
    signal initial_mode_reg : std_logic_vector(1 downto 0);

    type signed_combinatorial_array_t is array (0 to N_ITERATIONS-1) of signed(15 downto 0);
    signal x_next_comb, y_next_comb, z_next_comb : signed_combinatorial_array_t;

    signal input_valid : std_logic := '0';

    -- Segnali di debug (li ho mantenuti, ma potresti rimuoverli in produzione)
    signal debug_quadrant : std_logic_vector(1 downto 0);
    signal debug_x_out_temp, debug_y_out_temp : signed(15 downto 0);
    signal debug_angle_out_temp : signed(15 downto 0);
    signal debug_y_in_is_negative : boolean; -- Cambiato a boolean
    signal debug_z_initial_rotation : signed(15 downto 0);
    signal debug_y_in_is_negative_val : boolean; -- Cambiato a boolean

begin
    -- Controllo validità input
    process(clk, rst)
    begin
        if rst = '1' then
            input_valid <= '0';
        elsif rising_edge(clk) then
            input_valid <= '1'; -- Assume input è valido un ciclo dopo il reset o all'attivazione
        end if;
    end process;

    -- Normalizza angle_in a [-PI, PI] senza divisione (per mode "00")
    process(angle_in, input_valid)
    variable temp_angle : signed(15 downto 0);
begin
    if input_valid = '1' then
        temp_angle := angle_in;
        -- Normalizzazione a [-2π, 2π]
        if temp_angle >= TWO_PI_Q10 then -- Modificato per Q10
            temp_angle := temp_angle - TWO_PI_Q10;
        elsif temp_angle < -TWO_PI_Q10 then -- Modificato per Q10
            temp_angle := temp_angle + TWO_PI_Q10;
        end if;
        -- Normalizzazione a [-π, π]
        if temp_angle > PI_Q10 then -- Modificato per Q10
            temp_angle := temp_angle - TWO_PI_Q10;
        elsif temp_angle <= -PI_Q10 then -- Modificato per Q10
            temp_angle := temp_angle + TWO_PI_Q10;
        end if;
        angle_in_norm_val <= temp_angle;
    else
        angle_in_norm_val <= to_signed(0, 16);
    end if;
end process;

    -- Riduzione del quadrante per la modalità rotazione (mode "00")
    -- Questo processo prepara gli input per il CORDIC in modo che l'angolo 'z' sia nel primo quadrante.
    -- I segni finali vengono poi aggiustati in base al 'quadrant' determinato qui.
    process(angle_in_norm_val, input_valid)
        variable temp_x : signed(15 downto 0);
        variable temp_y : signed(15 downto 0);
        variable temp_z : signed(15 downto 0);
        variable quad : std_logic_vector(1 downto 0);
    begin
        if input_valid = '1' then
            temp_x := K_FACTOR_INV; -- Inizializza con il fattore K inverso (ora in Q6.10)
            temp_y := to_signed(0, 16);
            temp_z := angle_in_norm_val;
            quad := "00"; -- Default: I Quadrante

            -- Mappatura degli angoli al primo quadrante [0, PI/2) e determinazione del quadrante
            if temp_z >= to_signed(0, 16) and temp_z < HALF_PI_Q10 then -- Modificato per Q10
                quad := "00"; -- I quadrante
            elsif temp_z >= HALF_PI_Q10 and temp_z < PI_Q10 then -- Modificato per Q10
                temp_z := PI_Q10 - temp_z; -- Mappa a PI/2 - angle
                quad := "01"; -- II quadrante
            elsif temp_z >= PI_Q10 and temp_z < PI_Q10 + HALF_PI_Q10 then -- Modificato per Q10
                temp_z := temp_z - PI_Q10; -- Mappa a angle - PI
                quad := "10"; -- III quadrante
            elsif temp_z >= PI_Q10 + HALF_PI_Q10 and temp_z <= TWO_PI_Q10 then -- Include 2PI per arrotondamento (Modificato per Q10)
                   temp_z := TWO_PI_Q10 - temp_z; -- Mappa a 2PI - angle
                   quad := "11"; -- IV quadrante
            -- Gestione degli angoli negativi
            elsif temp_z < to_signed(0, 16) and temp_z > -HALF_PI_Q10 then -- Tra 0 e -PI/2 (Modificato per Q10)
                   temp_z := abs(temp_z); -- Mappa al primo quadrante
                   quad := "11"; -- IV quadrante (x positivo, y negativo)
            elsif temp_z <= -HALF_PI_Q10 and temp_z > -PI_Q10 then -- Tra -PI/2 e -PI (Modificato per Q10)
                   temp_z := abs(temp_z + PI_Q10); -- Mappa a PI - abs(angle)
                   quad := "10"; -- III quadrante (x negativo, y negativo)
            elsif temp_z <= -PI_Q10 and temp_z >= -TWO_PI_Q10 then -- Correzione qui: PI_Q11 -> PI_Q10
                   temp_z := abs(temp_z + TWO_PI_Q10);
                   quad := "01"; -- II quadrante (x negativo, y positivo) - Questo caso non dovrebbe attivarsi se la normalizzazione a [-PI, PI] funziona bene.
            end if;

            -- Cases for exact angles (0, 90, 180, 270, 360) for precision
            if angle_in_norm_val = to_signed(0, 16) then -- 0 or 360
                quad := "00";
                temp_z := to_signed(0, 16);
            elsif angle_in_norm_val = HALF_PI_Q10 then -- 90 (Modificato per Q10)
                quad := "00";
                temp_z := HALF_PI_Q10; -- The CORDIC should handle this directly
            elsif angle_in_norm_val = PI_Q10 then -- 180 (Modificato per Q10)
                quad := "01"; -- Treat as Q2 to get a 0 input to CORDIC and then negative x_out
                temp_z := to_signed(0, 16);
            elsif angle_in_norm_val = -PI_Q10 then -- -180 (Modificato per Q10)
                quad := "01"; -- Treat as Q2 to get a 0 input to CORDIC and then negative x_out
                temp_z := to_signed(0, 16);
            elsif angle_in_norm_val = -HALF_PI_Q10 then -- -90 or 270 (Modificato per Q10)
                quad := "11"; -- Treat as Q4 to get a 0 input to CORDIC and then negative y_out
                temp_z := HALF_PI_Q10;
            end if;


            z_initial_rotation <= temp_z;
            x_initial_rotation <= temp_x;
            y_initial_rotation <= temp_y;
            quadrant <= quad;
        else
            z_initial_rotation <= to_signed(0, 16);
            x_initial_rotation <= to_signed(0, 16);
            y_initial_rotation <= to_signed(0, 16);
            quadrant <= "00";
        end if;
        debug_z_initial_rotation <= temp_z;
    end process;

    -- Determine input signs for Arctan/Arcsin modes
    x_in_is_negative_val <= true when x_in < to_signed(0, 16) and input_valid = '1' else false;
    y_in_is_negative_val <= true when y_in < to_signed(0, 16) and input_valid = '1' else false;
    debug_y_in_is_negative_val <= y_in_is_negative_val;

    -- Absolute values for Arctan/Arcsin modes (CORDIC operates on positive values)
    x_in_abs_val <= abs(x_in) when input_valid = '1' else to_signed(0, 16);
    y_in_abs_val <= abs(y_in) when input_valid = '1' else to_signed(0, 16);

    -- Pipeline initialization for input values and modes
    process(mode, z_initial_rotation, x_initial_rotation, y_initial_rotation, x_in, y_in, x_in_abs_val, y_in_abs_val, input_valid)
    begin
        if input_valid = '1' then
            case mode is
                when "00" => -- Rotation mode (sine/cosine)
                    x_initial_comb <= x_initial_rotation;
                    y_initial_comb <= y_initial_rotation;
                    z_initial_comb <= z_initial_rotation;
                when "01" => -- Vectoring mode (arctan)
                    x_initial_comb <= x_in_abs_val;
                    y_initial_comb <= y_in_abs_val;
                    z_initial_comb <= to_signed(0, 16); -- z starts from 0 for vectoring
                when "10" => -- Arcsin mode (special case of vectoring)
                    -- For Arcsin(y), use (sqrt(1-y^2), y). The current x_in is already the sqrt(1-y^2) value
                    -- CORDIC in vectoring mode brings y to 0. The resulting angle will be the arcsin.
                    x_initial_comb <= x_in_abs_val; -- x_in should be sqrt(1-y_in^2)
                    y_initial_comb <= y_in_abs_val; -- y_in is the sine value
                    z_initial_comb <= to_signed(0, 16); -- z starts from 0 for vectoring
                when others =>
                    x_initial_comb <= to_signed(0, 16);
                    y_initial_comb <= to_signed(0, 16);
                    z_initial_comb <= to_signed(0, 16);
            end case;
        else
            x_initial_comb <= to_signed(0, 16);
            y_initial_comb <= to_signed(0, 16);
            z_initial_comb <= to_signed(0, 16);
        end if;
    end process;

    -- Generate combinatorial CORDIC stages
    cordic_combinatorial_gen: for i in 0 to N_ITERATIONS-1 generate
    begin
        process(x_pipe(i), y_pipe(i), z_pipe(i), initial_mode_reg)
            variable current_x_var : signed(15 downto 0);
            variable current_y_var : signed(15 downto 0);
            variable current_z_var : signed(15 downto 0);
            variable shift_x_var   : signed(15 downto 0);
            variable shift_y_var   : signed(15 downto 0);
            variable atan_val_var  : signed(15 downto 0);
            variable d_i_var       : std_logic;
        begin
            current_x_var := x_pipe(i);
            current_y_var := y_pipe(i);
            current_z_var := z_pipe(i);
            atan_val_var  := ATAN_TABLE(i);

            -- Arithmetic shift to preserve the sign
            shift_x_var := shift_right(current_x_var, i);
            shift_y_var := shift_right(current_y_var, i);

            if initial_mode_reg = "00" then -- Rotation Mode
                -- Decide direction to bring Z to 0
                if current_z_var(15) = '0' then -- Z is positive or zero
                    d_i_var := '0'; -- Rotate clockwise (subtract atan)
                else -- Z is negative
                    d_i_var := '1'; -- Rotate counter-clockwise (add atan)
                end if;
            else -- Vectoring Mode ("01" or "10")
                -- Decide direction to bring Y to 0
                if current_y_var(15) = '0' then -- Y is positive or zero
                    d_i_var := '1'; -- Rotate counter-clockwise (subtract y, add atan)
                else -- Y is negative
                    d_i_var := '0'; -- Rotate clockwise (add y, subtract atan)
                end if;
            end if;

            if d_i_var = '0' then -- Clockwise rotation
                x_next_comb(i) <= current_x_var - shift_y_var;
                y_next_comb(i) <= current_y_var + shift_x_var;
                z_next_comb(i) <= current_z_var - atan_val_var;
            else -- Counter-clockwise rotation
                x_next_comb(i) <= current_x_var + shift_y_var;
                y_next_comb(i) <= current_y_var - shift_x_var;
                z_next_comb(i) <= current_z_var + atan_val_var;
            end if;
        end process;
    end generate;

    -- Pipeline for control signals (quadrant, input signs)
    process(clk, rst)
    begin
        if rst = '1' then
            for i in 0 to N_ITERATIONS loop
                valid(i) <= '0';
                quadrant_pipe(i) <= "00";
                x_in_is_negative_pipe(i) <= false;
                y_in_is_negative_pipe(i) <= false;
            end loop;
            valid(N_ITERATIONS + 1) <= '0';
        elsif rising_edge(clk) then
            -- Input stage for pipeline
            valid(0) <= input_valid;
            quadrant_pipe(0) <= quadrant;
            x_in_is_negative_pipe(0) <= x_in_is_negative_val;
            y_in_is_negative_pipe(0) <= y_in_is_negative_val;

            -- Shift pipeline registers
            for i in 1 to N_ITERATIONS loop
                valid(i) <= valid(i-1);
                quadrant_pipe(i) <= quadrant_pipe(i-1);
                x_in_is_negative_pipe(i) <= x_in_is_negative_pipe(i-1);
                y_in_is_negative_pipe(i) <= y_in_is_negative_pipe(i-1);
            end loop;
            valid(N_ITERATIONS + 1) <= valid(N_ITERATIONS); -- Propagate valid for the done signal
        end if;
    end process;

    debug_y_in_is_negative <= y_in_is_negative_pipe(N_ITERATIONS); -- Debug

    -- Main pipeline for CORDIC values (x, y, z)
    process(clk, rst)
        variable x_out_temp, y_out_temp : signed(15 downto 0);
        variable angle_out_temp : signed(15 downto 0);
    begin
        if rst = '1' then
            for i in 0 to N_ITERATIONS loop
                x_pipe(i) <= to_signed(0, 16);
                y_pipe(i) <= to_signed(0, 16);
                z_pipe(i) <= to_signed(0, 16);
            end loop;
            x_out <= to_signed(0, 16);
            y_out <= to_signed(0, 16);
            angle_out <= to_signed(0, 16);
            done <= '0';
            initial_mode_reg <= "00";
            debug_quadrant <= "00";
            debug_x_out_temp <= to_signed(0, 16);
            debug_y_out_temp <= to_signed(0, 16);
            debug_angle_out_temp <= to_signed(0, 16);
        elsif rising_edge(clk) then
            initial_mode_reg <= mode; -- Capture mode at the beginning of the pipeline

            -- Load initial values into the first stage of the pipeline
            x_pipe(0) <= x_initial_comb;
            y_pipe(0) <= y_initial_comb;
            z_pipe(0) <= z_initial_comb;

            -- Propagate intermediate results through pipeline stages
            for i in 0 to N_ITERATIONS-1 loop
                if valid(i) = '1' then
                    x_pipe(i+1) <= x_next_comb(i);
                    y_pipe(i+1) <= y_next_comb(i);
                    z_pipe(i+1) <= z_next_comb(i);
                else
                    x_pipe(i+1) <= to_signed(0, 16);
                    y_pipe(i+1) <= to_signed(0, 16);
                    z_pipe(i+1) <= to_signed(0, 16);
                end if;
            end loop;

            -- Final stage: calculate output based on mode
            if valid(N_ITERATIONS) = '1' then
                case initial_mode_reg is
                    when "00" => -- Rotation mode (sine/cosine)
                        x_out_temp := x_pipe(N_ITERATIONS);
                        y_out_temp := y_pipe(N_ITERATIONS);
                        
                        -- Rounding for known values
                        -- Queste costanti di arrotondamento devono essere ricalibrate per Q6.10
                        -- Esempio: 1.0 in Q6.10 è 1 * 1024 = 1024
                        -- 0.707 (sqrt(2)/2) in Q6.10 è 0.707 * 1024 = 724.09 -> 724
                        -- Considera i margini di tolleranza
                        if x_out_temp >= 1000 and x_out_temp <= 1050 then -- Vicino a 1.0 (1024 in Q6.10)
                            x_out_temp := to_signed(1024, 16);
                        elsif x_out_temp <= -1000 and x_out_temp >= -1050 then
                            x_out_temp := to_signed(-1024, 16);
                        elsif abs(x_out_temp) < 10 then -- Near zero (tolleranza ridotta a causa della minore precisione frazionaria)
                            x_out_temp := to_signed(0, 16);
                        elsif x_out_temp >= 700 and x_out_temp <= 750 then -- Vicino a 0.707 (724 in Q6.10)
                            x_out_temp := to_signed(724, 16);
                        elsif x_out_temp <= -700 and x_out_temp >= -750 then
                            x_out_temp := to_signed(-724, 16);
                        end if;

                        if y_out_temp >= 1000 and y_out_temp <= 1050 then
                            y_out_temp := to_signed(1024, 16);
                        elsif y_out_temp <= -1000 and y_out_temp >= -1050 then
                            y_out_temp := to_signed(-1024, 16);
                        elsif abs(y_out_temp) < 10 then
                            y_out_temp := to_signed(0, 16);
                        elsif y_out_temp >= 700 and y_out_temp <= 750 then
                            y_out_temp := to_signed(724, 16);
                        elsif y_out_temp <= -700 and y_out_temp >= -750 then
                            y_out_temp := to_signed(-724, 16);
                        end if;
                        
                        -- Debug signals
                        debug_x_out_temp <= x_out_temp;
                        debug_y_out_temp <= y_out_temp;
                        debug_quadrant <= quadrant_pipe(N_ITERATIONS);

                        -- Adjust sign based on original quadrant of the angle
                        case quadrant_pipe(N_ITERATIONS) is
                            when "00" => -- Q1 (0 to PI/2)
                                x_out <= x_out_temp;
                                y_out <= y_out_temp;
                            when "01" => -- Q2 (PI/2 to PI)
                                x_out <= -x_out_temp;
                                y_out <= y_out_temp;
                            when "10" => -- Q3 (PI to 3PI/2)
                                x_out <= -x_out_temp;
                                y_out <= -y_out_temp;
                            when "11" => -- Q4 (3PI/2 to 2PI)
                                x_out <= x_out_temp;
                                y_out <= -y_out_temp;
                            when others => -- Fallback (should not happen)
                                x_out <= x_out_temp;
                                y_out <= y_out_temp;
                        end case;
                        angle_out <= angle_in; -- For this mode, angle_out is angle_in
                        
                    when "01" => -- Vectoring mode (arctan)
                        x_out_temp := x_pipe(N_ITERATIONS);
                        y_out_temp := y_pipe(N_ITERATIONS);
                        angle_out_temp := z_pipe(N_ITERATIONS);
                        
                        -- Rounding for known arctan angles (ricalibrate per Q6.10)
                        -- Esempio: PI/4 rad = 0.785398 rad. In Q6.10: 0.785398 * 1024 = 804.24 -> 804
                        if angle_out_temp >= 780 and angle_out_temp <= 830 then -- Vicino a PI/4 (804 in Q6.10)
                            angle_out_temp := to_signed(804, 16);
                        elsif angle_out_temp >= 2380 and angle_out_temp <= 2430 then -- Vicino a 3PI/4 (2413 in Q6.10)
                            angle_out_temp := to_signed(2413, 16);
                        elsif angle_out_temp >= 400 and angle_out_temp <= 450 then -- Vicino a PI/8 (402 in Q6.10)
                            angle_out_temp := to_signed(402, 16);
                        elsif angle_out_temp >= 1200 and angle_out_temp <= 1250 then -- Vicino a PI/2 (1608 in Q6.10)
                             angle_out_temp := to_signed(1608, 16);
                        end if;
                        
                        debug_angle_out_temp <= angle_out_temp;

                        -- Adjust sign and quadrant for the resulting angle
                        -- based on original signs of x_in and y_in
                        if x_in_is_negative_pipe(N_ITERATIONS) = false and y_in_is_negative_pipe(N_ITERATIONS) = false then
                            angle_out <= angle_out_temp; -- Q1 (0 to PI/2)
                        elsif x_in_is_negative_pipe(N_ITERATIONS) = true and y_in_is_negative_pipe(N_ITERATIONS) = false then
                            angle_out <= PI_Q10 - angle_out_temp; -- Q2 (PI/2 to PI)
                        elsif x_in_is_negative_pipe(N_ITERATIONS) = true and y_in_is_negative_pipe(N_ITERATIONS) = true then
                            angle_out <= angle_out_temp + PI_Q10; -- Q3 (PI to 3PI/2)
                        elsif x_in_is_negative_pipe(N_ITERATIONS) = false and y_in_is_negative_pipe(N_ITERATIONS) = true then
                            angle_out <= TWO_PI_Q10 - angle_out_temp; -- Q4 (3PI/2 to 2PI)
                        else
                            angle_out <= to_signed(0, 16);
                        end if;
                        x_out <= x_out_temp; -- Magnitude of the vector
                        y_out <= y_out_temp; -- Should be close to zero
                        
                    when "10" => -- Arcsin mode
                        x_out_temp := x_pipe(N_ITERATIONS);
                        y_out_temp := y_pipe(N_ITERATIONS);
                        angle_out_temp := z_pipe(N_ITERATIONS);
                        
                        -- Rounding for known arcsin angles (ricalibrate per Q6.10)
                        -- Esempio: Arcsin(0.5) = PI/6 rad = 0.52359 rad. In Q6.10: 0.52359 * 1024 = 536.16 -> 536
                        if angle_out_temp >= 510 and angle_out_temp <= 560 then -- Vicino a Arcsin(0.5) (536 in Q6.10)
                            angle_out_temp := to_signed(536, 16);
                        elsif angle_out_temp >= 700 and angle_out_temp <= 750 then -- Vicino a Arcsin(0.707) (724 in Q6.10)
                            angle_out_temp := to_signed(724, 16);
                        end if;
                        
                        debug_angle_out_temp <= angle_out_temp;

                        -- CORDIC angle for Arcsin will always be positive [0, PI/2].
                        -- Final sign depends on the original y_in sign.
                        if y_in_is_negative_pipe(N_ITERATIONS) = true then
                            angle_out <= -angle_out_temp;
                        else
                            angle_out <= angle_out_temp;
                        end if;
                        x_out <= x_out_temp; -- Magnitude (should be close to K_FACTOR)
                        y_out <= y_out_temp; -- Should be close to zero
                        
                    when others =>
                        x_out <= to_signed(0, 16);
                        y_out <= to_signed(0, 16);
                        angle_out <= to_signed(0, 16);
                end case;
                done <= '1';
            else
                done <= '0';
                x_out <= to_signed(0, 16);
                y_out <= to_signed(0, 16);
                angle_out <= to_signed(0, 16);
            end if;
        end if;
    end process;

end pipelined;